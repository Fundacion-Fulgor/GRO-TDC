** sch_path: /home/designer/shared/GRO-TDC/std_cells/XOR.sch
.subckt XOR OUT A VDD B VSS
*.PININFO VDD:B VSS:B A:I B:I OUT:O
x2 VDD net3 net2 B VSS AND
x4 VDD net3 A VSS INV_D1
x5 VDD net1 B VSS INV_D1
x1 VDD OUT net2 net4 VSS OR
x3 VDD A net4 net1 VSS AND
.ends

* expanding   symbol:  /home/designer/shared/GRO-TDC/std_cells/AND.sym # of pins=5
** sym_path: /home/designer/shared/GRO-TDC/std_cells/AND.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/AND.sch
.subckt AND VDD VA VOUT VB VSS
*.PININFO VDD:B VSS:B VA:I VB:I VOUT:O
x1 VDD VA net1 VB VSS NAND
x2 VDD VOUT net1 VSS INV_D1
.ends


* expanding   symbol:  /home/designer/shared/GRO-TDC/std_cells/INV_D1.sym # of pins=4
** sym_path: /home/designer/shared/GRO-TDC/std_cells/INV_D1.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/INV_D1.sch
.subckt INV_D1 VDD VOUT VIN VSS
*.PININFO VDD:B VSS:B VOUT:O VIN:I
M2 VOUT VIN VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/designer/shared/GRO-TDC/std_cells/OR.sym # of pins=5
** sym_path: /home/designer/shared/GRO-TDC/std_cells/OR.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/OR.sch
.subckt OR VDD VOUT VA VB VSS
*.PININFO VDD:B VSS:B VA:I VB:I VOUT:O
x2 VDD VOUT net1 VSS INV_D1
x1 VDD net1 VA VB VSS NOR
.ends


* expanding   symbol:  /home/designer/shared/GRO-TDC/std_cells/NAND.sym # of pins=5
** sym_path: /home/designer/shared/GRO-TDC/std_cells/NAND.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/NAND.sch
.subckt NAND VDD VA VOUT VB VSS
*.PININFO VDD:B VSS:B VA:I VB:I VOUT:O
M1 net1 VB VSS VSS sg13_lv_nmos w=0.45u l=0.13u ng=1 m=1
M2 VOUT VA net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M3 VOUT VB VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M4 VOUT VA VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/designer/shared/GRO-TDC/std_cells/NOR.sym # of pins=5
** sym_path: /home/designer/shared/GRO-TDC/std_cells/NOR.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/NOR.sch
.subckt NOR VDD VOUT VA VB VSS
*.PININFO VDD:B VSS:B VA:I VB:I VOUT:O
M1 VOUT VA VSS VSS sg13_lv_nmos w=0.45u l=0.13u ng=1 m=1
M2 VOUT VB VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M3 VOUT VB net1 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M4 net1 VA VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends

