** sch_path: /home/designer/shared/GRO-TDC/std_cells/NOR.sch
.subckt NOR VDD VOUT VA VB VSS
*.PININFO VDD:B VSS:B VA:I VB:I VOUT:O
M1 VOUT VA VSS VSS sg13_lv_nmos w=0.45u l=0.13u ng=1 m=1
M2 VOUT VB VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M3 VOUT VB net1 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M4 net1 VA VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends
