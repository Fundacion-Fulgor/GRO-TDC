* Extracted by KLayout with SG13G2 LVS runset on : 25/01/2026 23:58

.SUBCKT NOR VB
M$1 \$3 VB \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 \$1 \$5 \$3 \$1 sg13_lv_nmos L=0.13u W=0.45u AS=0.153p AD=0.153p PS=1.58u
+ PD=1.58u
M$3 \$2 \$5 \$6 \$2 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$4 \$6 VB \$3 \$2 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS NOR
