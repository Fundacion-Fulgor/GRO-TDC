* Extracted by KLayout with SG13G2 LVS runset on : 23/01/2026 18:55

.SUBCKT NAND_D2
M$1 \$5 \$4 \$6 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
M$2 \$6 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.9u AS=0.306p AD=0.306p PS=2.48u
+ PD=2.48u
M$3 \$5 \$3 \$2 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
M$4 \$2 \$4 \$5 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS NAND_D2
