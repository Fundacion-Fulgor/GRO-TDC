** sch_path: /foss/designs/GRO-TDC/std_cells/MUX_8_1.sch
**.subckt MUX_8_1 VINA VINB VDD VOUT CTRL[2],CTRL[1],CTRL[0] VINC VSS VIND
*.iopin VSS
*.opin VOUT
*.iopin VDD
*.ipin VINA
*.ipin VINB
*.ipin VINC
*.ipin VIND
*.ipin VS[2],VS[1],VS[0]
*.ipin VINE
*.ipin VINF
*.ipin VING
*.ipin VINH
x7 VDD net1 VOUT VS[2] net2 VSS MUX_2_1
x8 VINA VINB VDD net1 VS[1] VS[0] VINC VSS VIND VS[1] MUX_4_1
x9 VINE VINF VDD net2 VS[1] VS[0] VING VSS VINH VS[1] MUX_4_1
**.ends

* expanding   symbol:  /foss/designs/PhaseInterpolator/Custom_std_cells/MUX_2_1.sym # of pins=6
** sym_path: /foss/designs/PhaseInterpolator/Custom_std_cells/MUX_2_1.sym
** sch_path: /foss/designs/PhaseInterpolator/Custom_std_cells/MUX_2_1.sch
.subckt MUX_2_1 VDD VINA VOUT VS VINB VSS
*.opin VOUT
*.ipin VINA
*.ipin VINB
*.ipin VS
*.iopin VDD
*.iopin VSS
x1 VOUT net1 VS net2 VDD VSS tg_custom
x2 VOUT VS net1 net3 VDD VSS tg_custom
x3 VDD net1 VS VSS inv
x4 VDD net2 VINA VSS inv_PI
x5 VDD net3 VINB VSS inv_PI
x6[3] VOUT VSS VDD net2 VDD VSS tg_custom
x6[2] VOUT VSS VDD net2 VDD VSS tg_custom
x6[1] VOUT VSS VDD net2 VDD VSS tg_custom
x6[0] VOUT VSS VDD net2 VDD VSS tg_custom
x7[3] VOUT VSS VDD net3 VDD VSS tg_custom
x7[2] VOUT VSS VDD net3 VDD VSS tg_custom
x7[1] VOUT VSS VDD net3 VDD VSS tg_custom
x7[0] VOUT VSS VDD net3 VDD VSS tg_custom
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/MUX_4_1.sym # of pins=9
** sym_path: /foss/designs/GRO-TDC/std_cells/MUX_4_1.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/MUX_4_1.sch
.subckt MUX_4_1 VINA VINB VDD VOUT VS[1] VS[0] VINC VSS VIND VST
*.opin VOUT
*.iopin VDD
*.iopin VSS
*.ipin VINA
*.ipin VINB
*.ipin VINC
*.ipin VIND
*.ipin VS[1],VS[0]
*.ipin VST
x3 VDD VINC net2 VS[1] VIND VSS MUX_2_1
x4 VDD VINA net1 VS[0] VINB VSS MUX_2_1
x5 VDD net1 VOUT VST net2 VSS MUX_2_1
.ends


* expanding   symbol:  /foss/designs/PhaseInterpolator/Custom_std_cells/tg_custom.sym # of pins=6
** sym_path: /foss/designs/PhaseInterpolator/Custom_std_cells/tg_custom.sym
** sch_path: /foss/designs/PhaseInterpolator/Custom_std_cells/tg_custom.sch
.subckt tg_custom VOUT VSN VSP VIN VBP VBN
*.iopin VIN
*.iopin VSN
*.iopin VOUT
*.iopin VSP
*.iopin VBN
*.iopin VBP
XM1 VOUT VSN VIN VBN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 VOUT VSP VIN VBP sg13_lv_pmos w=0.3u l=0.13u ng=2 m=1
.ends


* expanding   symbol:  /foss/designs/PhaseInterpolator/Custom_std_cells/inv.sym # of pins=4
** sym_path: /foss/designs/PhaseInterpolator/Custom_std_cells/inv.sym
** sch_path: /foss/designs/PhaseInterpolator/Custom_std_cells/inv.sch
.subckt inv VDD VOUT VIN VSS
*.iopin VDD
*.iopin VSS
*.opin VOUT
*.ipin VIN
XM2 VOUT VIN VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/PhaseInterpolator/Custom_std_cells/inv_PI.sym # of pins=4
** sym_path: /foss/designs/PhaseInterpolator/Custom_std_cells/inv_PI.sym
** sch_path: /foss/designs/PhaseInterpolator/Custom_std_cells/inv_PI.sch
.subckt inv_PI VDD VOUT VIN VSS
*.iopin VDD
*.iopin VSS
*.opin VOUT
*.ipin VIN
XM2 VOUT VIN VDD VDD sg13_lv_pmos w=0.45u l=0.13u ng=3 m=1
XM1 VOUT VIN VSS VSS sg13_lv_nmos w=0.3u l=0.13u ng=2 m=1
.ends

.end
