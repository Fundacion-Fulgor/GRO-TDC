* Extracted by KLayout with SG13G2 LVS runset on : 21/01/2026 22:49

.SUBCKT INV3
X$4 \$4 \$5 \$2 \$3 INV_D1
X$5 \$4 \$5 \$2 \$3 INV_D1
X$6 \$4 \$5 \$2 \$3 INV_D1
X$7 \$4 \$5 \$2 \$3 INV_D1
X$8 \$4 \$5 \$I3 \$1 INV_D1
X$9 \$4 \$5 \$1 \$2 INV_D1
X$10 \$4 \$5 \$1 \$2 INV_D1
.ENDS INV3

.SUBCKT INV_D1 \$1 \$2 \$3 \$4
M$1 \$2 \$3 \$4 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
M$2 \$1 \$3 \$4 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS INV_D1
