* Extracted by KLayout with SG13G2 LVS runset on : 25/01/2026 21:46

.SUBCKT INV_D2
M$1 \$1 \$4 \$3 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
M$2 \$2 \$4 \$3 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS INV_D2
