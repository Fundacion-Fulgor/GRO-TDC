* Extracted by KLayout with SG13G2 LVS runset on : 25/01/2026 23:34

.SUBCKT Modi_Buffers VDD IN0|IN2 IN0 K0 K1 K2 IN0$1 VSS IN0$2 IN0|IN1 IN0$3
M$1 IN0$1 K0 \$11 VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$2 \$11 K0 VSS VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$3 IN0|IN2 K1 \$12 VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$4 \$12 K1 VSS VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$5 IN0 K2 \$13 VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$6 \$13 K2 VSS VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$7 VSS IN0$2 IN0$1 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p
+ PS=2.68u PD=2.68u
M$8 VSS IN0$1 K0 VSS sg13_lv_nmos L=0.13u W=0.6u AS=0.204p AD=0.204p PS=2.56u
+ PD=2.56u
M$9 VSS IN0|IN1 IN0|IN2 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p
+ PS=2.68u PD=2.68u
M$10 VSS IN0|IN2 K1 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p
+ PS=2.68u PD=2.68u
M$11 VSS IN0$3 IN0 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p PS=2.68u
+ PD=2.68u
M$12 VSS IN0 K2 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p PS=2.68u
+ PD=2.68u
M$19 IN0$1 K0 VDD VDD sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$20 IN0|IN2 K1 VDD VDD sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$21 IN0 K2 VDD VDD sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$22 VDD IN0$2 IN0$1 VDD sg13_lv_pmos L=0.13u W=0.6u AS=0.204p AD=0.204p
+ PS=2.56u PD=2.56u
M$23 VDD IN0$1 K0 VDD sg13_lv_pmos L=0.13u W=0.6u AS=0.204p AD=0.204p PS=2.56u
+ PD=2.56u
M$24 VDD IN0|IN1 IN0|IN2 VDD sg13_lv_pmos L=0.13u W=0.6u AS=0.204p AD=0.204p
+ PS=2.56u PD=2.56u
M$25 VDD IN0|IN2 K1 VDD sg13_lv_pmos L=0.13u W=0.6u AS=0.204p AD=0.204p
+ PS=2.56u PD=2.56u
M$26 VDD IN0$3 IN0 VDD sg13_lv_pmos L=0.13u W=0.6u AS=0.204p AD=0.204p PS=2.56u
+ PD=2.56u
M$27 VDD IN0 K2 VDD sg13_lv_pmos L=0.13u W=0.6u AS=0.204p AD=0.204p PS=2.56u
+ PD=2.56u
.ENDS Modi_Buffers
