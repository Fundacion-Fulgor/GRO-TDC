* Extracted by KLayout with SG13G2 LVS runset on : 07/01/2026 20:41

.SUBCKT INV_D1 VSS VDD VOUT VIN
M$1 VSS VIN VOUT VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$2 VDD VIN VOUT VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS INV_D1
