** sch_path: /home/designer/shared/GRO-TDC/std_cells/TG_2C.sch
.subckt TG_2C VCTRLN VSS VOUT VIN VDD VCTRLP
*.PININFO VCTRLN:B VCTRLP:B VOUT:O VIN:I VSS:B VDD:B
M1 VOUT VCTRLN VIN VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M2 VOUT VCTRLP VIN VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=2
.ends
