* Extracted by KLayout with SG13G2 LVS runset on : 28/01/2026 00:30

.SUBCKT GRO
X$4 \$8 \$3 \$1 \$7 INV3
X$5 \$7 \$3 \$1 \$2 INV3
X$77 \$2 \$3 \$1 \$8 INV3
X$81 \$1 \$12 \$11 \$20 INV_D1
X$82 \$1 \$12 \$11 \$20 INV_D1
X$83 \$1 \$12 \$11 \$20 INV_D1
X$84 \$1 \$12 \$11 \$20 INV_D1
X$85 \$1 \$12 \$20 \$16 INV_D1
X$86 \$1 \$12 \$20 \$16 INV_D1
X$87 \$1 \$12 \$20 \$16 INV_D1
X$88 \$1 \$12 \$20 \$16 INV_D1
X$89 \$1 \$12 \$20 \$16 INV_D1
X$90 \$1 \$12 \$20 \$16 INV_D1
X$91 \$1 \$12 \$20 \$16 INV_D1
X$92 \$1 \$12 \$20 \$16 INV_D1
X$93 \$1 \$12 \$16 \$9 INV_D1
X$94 \$1 \$12 \$16 \$9 INV_D1
X$95 \$1 \$12 \$16 \$9 INV_D1
X$96 \$1 \$12 \$16 \$9 INV_D1
X$97 \$1 \$12 \$16 \$9 INV_D1
X$98 \$1 \$12 \$16 \$9 INV_D1
X$99 \$1 \$12 \$16 \$9 INV_D1
X$100 \$1 \$12 \$16 \$9 INV_D1
X$101 \$1 \$12 \$16 \$9 INV_D1
X$102 \$1 \$12 \$16 \$9 INV_D1
X$103 \$1 \$12 \$16 \$9 INV_D1
X$104 \$1 \$12 \$16 \$9 INV_D1
X$105 \$1 \$12 \$16 \$9 INV_D1
X$106 \$1 \$12 \$16 \$9 INV_D1
X$107 \$1 \$12 \$16 \$9 INV_D1
X$108 \$1 \$12 \$16 \$9 INV_D1
X$109 \$1 \$12 \$23 \$11 INV_D1
X$112 \$1 \$12 \$23 \$11 INV_D1
M$1 \$12 \$11 \$7 \$12 sg13_lv_pmos L=0.13u W=4.8u AS=1.956p AD=1.956p
+ PS=26.08u PD=26.08u
M$33 \$3 \$9 \$12 \$12 sg13_lv_pmos L=0.13u W=4.8u AS=1.956p AD=1.956p
+ PS=26.08u PD=26.08u
M$65 \$1 \$9 \$2 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$66 \$1 \$9 \$3 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
.ENDS GRO

.SUBCKT INV3 \$3 \$4 \$5 \$I5
X$4 \$5 \$4 \$2 \$3 INV_D1
X$5 \$5 \$4 \$2 \$3 INV_D1
X$6 \$5 \$4 \$2 \$3 INV_D1
X$7 \$5 \$4 \$2 \$3 INV_D1
X$8 \$5 \$4 \$I5 \$1 INV_D1
X$9 \$5 \$4 \$1 \$2 INV_D1
X$10 \$5 \$4 \$1 \$2 INV_D1
.ENDS INV3

.SUBCKT INV_D1 \$1 \$2 \$3 \$4
M$1 \$2 \$3 \$4 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
M$2 \$1 \$3 \$4 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS INV_D1
