* Extracted by KLayout with SG13G2 LVS runset on : 25/01/2026 15:47

.SUBCKT SR_Latch VSS VS VR VDD QN QP
X$1 VR QN VDD VSS QP NOR
X$2 QP VS VDD VSS QN NOR
.ENDS SR_Latch

.SUBCKT NOR VB \$2 \$3 \$4 \$5
M$1 \$4 VB \$5 \$4 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 \$5 \$2 \$4 \$4 sg13_lv_nmos L=0.13u W=0.45u AS=0.153p AD=0.153p PS=1.58u
+ PD=1.58u
M$3 \$5 VB \$7 \$3 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$4 \$7 \$2 \$3 \$3 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS NOR
