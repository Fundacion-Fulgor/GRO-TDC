* Extracted by KLayout with SG13G2 LVS runset on : 24/01/2026 01:08

.SUBCKT FF_D_routed
X$1 \$3 \$1 VIA1_constraint
X$2 \$1 \$2 \$15 \$15 \$8 \$5 \$4 \$3 \$5 \$2 \$12 \$12 \$3 \$4 \$2 \$9 \$13
+ \$5 \$12 FF_D_placement
X$3 \$4 \$1 VIA1_constraint
X$4 \$13 \$1 VIA1_constraint
X$5 \$12 \$1 VIA1_constraint
X$6 \$12 \$1 VIA2_constraint
X$7 \$12 \$1 VIA3_constraint
X$8 \$12 \$1 VIA1_constraint
X$9 \$12 \$1 VIA3_constraint
X$10 \$12 \$1 VIA2_constraint
X$11 \$12 \$1 VIA1_constraint
X$12 \$12 \$1 VIA2_constraint
X$13 \$12 \$1 VIA2_constraint
X$14 \$2 \$1 VIA1_constraint
X$15 \$2 \$1 VIA2_constraint
X$16 \$5 \$1 VIA2_constraint
X$17 \$5 \$1 VIA1_constraint
X$18 \$2 \$1 VIA1_constraint
X$19 \$2 \$1 VIA2_constraint
X$20 \$2 \$1 VIA2_constraint
X$21 \$2 \$1 VIA2_constraint
X$22 \$5 \$1 VIA2_constraint
.ENDS FF_D_routed

.SUBCKT FF_D_placement \$1 \$I24 \$I23 \$I22 \$I21 \$I20 \$I19 \$I18 \$I17
+ \$I16 \$I15 \$I14 \$I13 \$I12 \$I11 \$I7 \$I6 \$I5 \$I4
X$1 \$1 \$I10 \$I7 \$I4 INV_D1
X$2 \$1 \$I20 \$I21 \$I7 \$I19 \$I24 \$I14 \$I13 HALF_B
X$3 \$1 \$I11 \$I7 \$I5 INV_D1
X$4 \$1 \$I22 \$I18 \$I16 \$I7 \$I17 \$I15 \$I23 HALF_A
X$5 \$1 \$I12 \$I7 \$I6 INV_D1
.ENDS FF_D_placement

.SUBCKT HALF_A \$1 \$2 \$3 \$5 \$10 \$13 \$I37 \$I18
X$1 \$1 \$11 \$10 \$2 INV_D1
X$2 \$5 \$13 \$I25 \$1 \$I18 \$4 TG_2C
X$3 \$13 \$5 \$I25 \$1 \$9 \$4 TG_2C
X$4 \$2 \$1 VIA1_constraint
X$5 \$1 \$3 \$10 \$9 INV_D1
X$6 \$13 \$1 VIA1_constraint
X$7 \$13 \$1 VIA2_constraint
X$8 \$13 \$1 VIA2_constraint
X$9 \$4 \$1 VIA1_constraint
X$10 \$I18 \$1 VIA1_constraint
X$11 \$4 \$1 VIA1_constraint
X$12 \$13 \$1 VIA1_constraint
X$13 \$9 \$1 VIA1_constraint
X$14 \$9 \$1 VIA1_constraint
X$15 \$4 \$1 VIA2_constraint
X$16 \$1 \$10 \$4 \$I37 \$3 NAND_D2
X$17 \$4 \$1 VIA2_constraint
X$18 \$4 \$1 VIA1_constraint
X$19 \$3 \$1 VIA1_constraint
.ENDS HALF_A

.SUBCKT HALF_B \$1 \$3 \$6 \$7 \$14 \$15 \$I52 \$I51
X$1 \$3 \$15 \$6 \$1 \$11 \$2 TG_2C
X$2 \$I52 \$2 \$6 \$1 \$14 NAND_D3
X$3 \$15 \$3 \$7 \$1 \$10 \$4 TG_2C
X$4 \$14 \$1 VIA2_constraint
X$5 \$14 \$1 VIA3_constraint
X$6 \$1 \$14 \$7 \$10 INV_D1
X$7 \$I51 \$1 \$11 \$6 INV_D3
X$8 \$10 \$1 VIA1_constraint
X$9 \$14 \$1 VIA1_constraint
X$10 \$14 \$1 VIA2_constraint
X$11 \$14 \$1 VIA3_constraint
X$12 \$15 \$1 VIA1_constraint
X$13 \$2 \$1 VIA1_constraint
X$14 \$11 \$1 VIA1_constraint
X$15 \$3 \$1 VIA1_constraint
X$16 \$3 \$1 VIA2_constraint
X$17 \$15 \$1 VIA2_constraint
X$18 \$3 \$1 VIA2_constraint
X$19 \$15 \$1 VIA1_constraint
X$20 \$4 \$1 VIA1_constraint
X$21 \$10 \$1 VIA1_constraint
X$22 \$3 \$1 VIA1_constraint
X$23 \$15 \$1 VIA2_constraint
.ENDS HALF_B

.SUBCKT NAND_D2 \$1 \$2 \$3 \$4 \$5
X$1 \$1 \$6 \$1 \$3 nmos$1
X$2 \$6 \$5 \$1 \$4 nmos$2
X$3 \$2 \$5 \$3 \$2 \$1 pmos$2
X$4 \$5 \$2 \$4 \$2 \$1 pmos$2
.ENDS NAND_D2

.SUBCKT VIA3_constraint \$1 \$2
.ENDS VIA3_constraint

.SUBCKT VIA2_constraint \$1 \$2
.ENDS VIA2_constraint

.SUBCKT VIA1_constraint \$1 \$2
.ENDS VIA1_constraint

.SUBCKT INV_D3 \$1 \$2 \$4 \$10
X$1 \$2 \$10 \$4 \$1 INV
X$2 \$2 \$10 \$4 \$1 INV
X$3 \$2 \$10 \$4 \$1 INV
M$1 \$4 \$1 \$2 \$2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$2 \$1 \$4 \$2 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$3 \$2 \$1 \$4 \$2 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$4 \$10 \$1 \$4 \$10 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$5 \$4 \$1 \$10 \$10 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$6 \$10 \$1 \$4 \$10 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$7 \$4 \$1 \$10 \$10 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$8 \$10 \$1 \$4 \$10 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.0555p
+ PS=0.74u PD=0.74u
M$9 \$4 \$1 \$10 \$10 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
.ENDS INV_D3

.SUBCKT TG_2C \$1 \$2 \$3 \$4 \$5 \$6
X$1 \$6 \$5 \$4 \$1 nmos
X$2 \$5 \$6 \$2 \$3 \$4 pmos
X$3 \$6 \$5 \$2 \$3 \$4 pmos
M$1 \$5 \$2 \$6 \$3 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$6 \$2 \$5 \$3 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
.ENDS TG_2C

.SUBCKT INV_D1 \$1 \$2 \$3 \$4
X$1 \$1 \$4 \$1 \$2 nmos$3
X$2 \$4 \$3 \$2 \$3 \$1 pmos$1
.ENDS INV_D1

.SUBCKT NAND_D3 \$1 \$2 \$3 \$4 \$5
X$1 \$3 \$5 \$1 \$3 \$4 pmos$3
X$2 \$5 \$6 \$4 \$1 nmos$4
X$3 \$6 \$4 \$4 \$2 nmos$1$1
X$4 \$5 \$3 \$2 \$3 \$4 pmos$3
.ENDS NAND_D3

.SUBCKT nmos$2 \$1 \$2 \$3 \$5
M$1 \$2 \$5 \$1 \$3 sg13_lv_nmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS nmos$2

.SUBCKT nmos$1 \$1 \$2 \$3 \$5
M$1 \$2 \$5 \$1 \$3 sg13_lv_nmos L=0.13u W=0.9u AS=0.306p AD=0.306p PS=2.48u
+ PD=2.48u
.ENDS nmos$1

.SUBCKT pmos$2 \$1 \$2 \$3 \$4 \$6
M$1 \$2 \$3 \$1 \$4 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS pmos$2

.SUBCKT INV \$1 \$2 \$3 \$4
X$1 \$1 \$3 \$1 \$4 nmos$5
X$2 \$3 \$2 \$4 \$2 \$1 pmos$4
X$3 \$2 \$3 \$4 \$2 \$1 pmos$4
.ENDS INV

.SUBCKT pmos \$1 \$2 \$3 \$4 \$6
.ENDS pmos

.SUBCKT nmos \$1 \$2 \$3 \$5
M$1 \$2 \$5 \$1 \$3 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS nmos

.SUBCKT pmos$1 \$1 \$2 \$3 \$4 \$6
M$1 \$2 \$3 \$1 \$4 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS pmos$1

.SUBCKT nmos$3 \$1 \$2 \$3 \$5
M$1 \$1 \$5 \$2 \$3 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS nmos$3

.SUBCKT nmos$4 \$1 \$2 \$3 \$5
M$1 \$1 \$5 \$2 \$3 sg13_lv_nmos L=0.13u W=0.45u AS=0.153p AD=0.153p PS=1.58u
+ PD=1.58u
.ENDS nmos$4

.SUBCKT nmos$1$1 \$1 \$2 \$3 \$5
M$1 \$1 \$5 \$2 \$3 sg13_lv_nmos L=0.13u W=1.35u AS=0.459p AD=0.459p PS=3.38u
+ PD=3.38u
.ENDS nmos$1$1

.SUBCKT pmos$3 \$1 \$2 \$3 \$4 \$6
M$1 \$1 \$3 \$2 \$4 sg13_lv_pmos L=0.13u W=0.45u AS=0.153p AD=0.153p PS=1.58u
+ PD=1.58u
.ENDS pmos$3

.SUBCKT pmos$4 \$1 \$2 \$3 \$4 \$6
.ENDS pmos$4

.SUBCKT nmos$5 \$1 \$2 \$3 \$5
.ENDS nmos$5
