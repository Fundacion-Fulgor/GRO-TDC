* Extracted by KLayout with SG13G2 LVS runset on : 25/01/2026 18:00

.SUBCKT INV05
M$1 \$1 \$5 \$3 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$3 \$5 \$4 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$3 \$2 \$5 \$4 \$2 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS INV05
