** sch_path: /home/designer/shared/GRO-TDC/std_cells/NAND_D2.sch
.subckt NAND_D2 VDD VA VOUT VB VSS
*.PININFO VDD:B VSS:B VA:I VB:I VOUT:O
M1 net1 VB VSS VSS sg13_lv_nmos w=0.9u l=0.13u ng=1 m=1
M2 VOUT VA net1 VSS sg13_lv_nmos w=0.3u l=0.13u ng=1 m=1
M3 VOUT VB VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M4 VOUT VA VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends
