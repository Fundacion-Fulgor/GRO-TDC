** sch_path: /foss/designs/GRO-TDC/GROTDC_SIM/tb_Counter_FA_6bits.sch
**.subckt tb_Counter_FA_6bits
V1 VSS GND 0
V3 B[0] VSS dc {B0}
V5 VDD VSS 1.2
V4 A[0] VSS dc {A0}
x1 S[5] S[4] S[3] S[2] S[1] S[0] A[5] A[4] A[3] A[2] A[1] A[0] VDD COUT B[5] B[4] B[3] B[2] B[1] B[0] VSS CIN Counter_FA_6bits
V2 A[1] VSS dc {A1}
V6 A[2] VSS dc {A2}
V7 A[3] VSS dc {A3}
V8 A[4] VSS dc {A4}
V9 A[5] VSS dc {A5}
V10 B[1] VSS dc {B1}
V11 B[2] VSS dc {B2}
V12 B[3] VSS dc {B3}
V13 B[4] VSS dc {B4}
V14 B[5] VSS dc {B5}
V15 CIN VSS dc {CI}
**** begin user architecture code



.param CI=0
.param A0=1
.param A1=1
.param A2=1
.param A3=1
.param A4=1
.param A5=1

.param B0=1
.param B1=1
.param B2=1
.param B3=1
.param B4=1
.param B5=1


.param temp=65
.control
save all
tran 500p 30n
*let sum0 = v(S[0])
*let sum1 = v(S[1])
*let sum2 = v(S[2])
*let sum3 = v(S[3])
*let sum4 = v(S[4])
*let sum5 = v(S[5])

*print sum0 sum1 sum2 sum3 sum4 sum5

write counter2_tb.raw
*set appendwrite
.endc




.lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/Counter_FA_6bits.sym # of pins=7
** sym_path: /foss/designs/GRO-TDC/std_cells/Counter_FA_6bits.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/Counter_FA_6bits.sch
.subckt Counter_FA_6bits S[5] S[4] S[3] S[2] S[1] S[0] A[5] A[4] A[3] A[2] A[1] A[0] VDD COUT B[5] B[4] B[3] B[2] B[1] B[0] VSS
+ CIN
*.iopin VDD
*.iopin VSS
*.ipin A[5],A[4],A[3],A[2],A[1],A[0]
*.ipin B[5],B[4],B[3],B[2],B[1],B[0]
*.ipin CIN
*.opin S[5],S[4],S[3],S[2],S[1],S[0]
*.opin COUT
x6 A[0] VDD B[0] S[0] VSS CIN net1 FA
x1 A[1] VDD B[1] S[1] VSS net1 net2 FA
x2 A[2] VDD B[2] S[2] VSS net2 net3 FA
x3 A[3] VDD B[3] S[3] VSS net3 net4 FA
x4 A[4] VDD B[4] S[4] VSS net4 net5 FA
x5 A[5] VDD B[5] S[5] VSS net5 COUT FA
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/FA.sym # of pins=7
** sym_path: /foss/designs/GRO-TDC/std_cells/FA.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/FA.sch
.subckt FA A VDD B S VSS CIN CSAL
*.ipin B
*.ipin A
*.ipin CIN
*.opin S
*.opin CSAL
*.iopin VDD
*.iopin VSS
x1 net2 B VDD CIN VSS XOR
x5 S A VDD net2 VSS XOR
x6 VDD net1 net4 net3 VSS OR
x7 VDD CSAL net1 net5 VSS OR
x2 VDD B net4 CIN VSS AND
x3 VDD B net3 A VSS AND
x4 VDD CIN net5 A VSS AND
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/XOR.sym # of pins=5
** sym_path: /foss/designs/GRO-TDC/std_cells/XOR.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/XOR.sch
.subckt XOR OUT A VDD B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
x2 VDD net3 net2 B VSS AND
x4 VDD net3 A VSS INV_D1
x5 VDD net1 B VSS INV_D1
x1 VDD OUT net2 net4 VSS OR
x3 VDD A net4 net1 VSS AND
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/OR.sym # of pins=5
** sym_path: /foss/designs/GRO-TDC/std_cells/OR.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/OR.sch
.subckt OR VDD VOUT VA VB VSS
*.iopin VDD
*.iopin VSS
*.ipin VA
*.ipin VB
*.opin VOUT
x2 VDD VOUT net1 VSS INV_D1
x1 VDD net1 VA VB VSS NOR
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/AND.sym # of pins=5
** sym_path: /foss/designs/GRO-TDC/std_cells/AND.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/AND.sch
.subckt AND VDD VA VOUT VB VSS
*.iopin VDD
*.iopin VSS
*.ipin VA
*.ipin VB
*.opin VOUT
x1 VDD VA net1 VB VSS NAND
x2 VDD VOUT net1 VSS INV_D1
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/INV_D1.sym # of pins=4
** sym_path: /foss/designs/GRO-TDC/std_cells/INV_D1.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/INV_D1.sch
.subckt INV_D1 VDD VOUT VIN VSS
*.iopin VDD
*.iopin VSS
*.opin VOUT
*.ipin VIN
XM2 VOUT VIN VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/NOR.sym # of pins=5
** sym_path: /foss/designs/GRO-TDC/std_cells/NOR.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/NOR.sch
.subckt NOR VDD VOUT VA VB VSS
*.iopin VDD
*.iopin VSS
*.ipin VA
*.ipin VB
*.opin VOUT
XM1 VOUT VA VSS VSS sg13_lv_nmos w=0.45u l=0.13u ng=1 m=1
XM2 VOUT VB VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM3 VOUT VB net1 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM4 net1 VA VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/NAND.sym # of pins=5
** sym_path: /foss/designs/GRO-TDC/std_cells/NAND.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/NAND.sch
.subckt NAND VDD VA VOUT VB VSS
*.iopin VDD
*.iopin VSS
*.ipin VA
*.ipin VB
*.opin VOUT
XM1 net1 VB VSS VSS sg13_lv_nmos w=0.45u l=0.13u ng=1 m=1
XM2 VOUT VA net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM3 VOUT VB VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM4 VOUT VA VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
