** sch_path: /home/designer/shared/GRO-TDC/std_cells/INV05.sch
.subckt INV05 VDD VOUT VIN VSS
*.PININFO VDD:B VSS:B VOUT:O VIN:I
M1 net1 VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M3 VOUT VIN VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M2 VOUT VIN net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends
