* Extracted by KLayout with SG13G2 LVS runset on : 24/01/2026 15:34

.SUBCKT TG_2C VOUT VIN
M$1 VIN \$2 VOUT \$3 sg13_lv_pmos L=0.13u W=0.3u AS=0.156p AD=0.156p PS=2.08u
+ PD=2.08u
M$3 VIN \$1 VOUT \$4 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
.ENDS TG_2C
