** sch_path: /home/designer/shared/GRO-TDC/std_cells/INV_D2.sch
.subckt INV_D2 VDD VOUT VIN VSS
*.PININFO VDD:B VSS:B VOUT:O VIN:I
M1 VOUT VIN VSS VSS sg13_lv_nmos w=0.3u l=0.13u ng=1 m=1
M2 VOUT VIN VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends
