** sch_path: /foss/designs/GRO-TDC/GROTDC_SIM/tb_TG_2C.sch
**.subckt tb_TG_2C
V1 VSS GND 0
V3 VIN1 VSS dc 0 ac 0 pulse(0, 1.2, 0, 1p, 1p, 10n, 20n)
V5 VDD VSS 1.2
x1 VCLK VSS VOUT VIN VDD VCLKN TG_2C
x10 VDD VCLK_N VCLK VSS INV_D1
V2 VCLK1 VSS dc 0 ac 0 pulse(0, 1.2, 3.5n, 10p, 10p, 5n, 10n)
x2 VDD net2 VOUT VSS INV_D1
x3 VDD VIN net1 VSS INV_D1
x4[2] VDD net1 VIN1 VSS INV_D1
x4[1] VDD net1 VIN1 VSS INV_D1
x4[0] VDD net1 VIN1 VSS INV_D1
x1[1] VDD VCLK VCLK1 VSS INV_D1
x1[0] VDD VCLK VCLK1 VSS INV_D1
R1 net2 VSS 1k m=1
**** begin user architecture code


.param temp=65
.control
save all
tran 50p 50n
*let clk0 = v(CLK)
*let VB0 = v(B0)


*plot VB0
*plot VB1
*plot clk0
*plot clk1

write counter_tb.raw
set appendwrite
.endc



.lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/TG_2C.sym # of pins=6
** sym_path: /foss/designs/GRO-TDC/std_cells/TG_2C.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/TG_2C.sch
.subckt TG_2C VCTRLN VSS VOUT VIN VDD VCTRLP
*.iopin VCTRLN
*.iopin VCTRLP
*.opin VOUT
*.ipin VIN
*.iopin VSS
*.iopin VDD
XM1 VOUT VCTRLN VIN VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 VOUT VCTRLP VIN VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=2
.ends


* expanding   symbol:  /foss/designs/GRO-TDC/std_cells/INV_D1.sym # of pins=4
** sym_path: /foss/designs/GRO-TDC/std_cells/INV_D1.sym
** sch_path: /foss/designs/GRO-TDC/std_cells/INV_D1.sch
.subckt INV_D1 VDD VOUT VIN VSS
*.iopin VDD
*.iopin VSS
*.opin VOUT
*.ipin VIN
XM2 VOUT VIN VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
XM1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
