** sch_path: /home/designer/shared/GRO-TDC/std_cells/INV3.sch
.subckt INV3 VDD VOUT VIN VSS
*.PININFO VDD:B VSS:B VOUT:O VIN:I
x2 VDD net2 VIN VSS INV_D1
x1[1] VDD net1 net2 VSS INV_D1
x1[0] VDD net1 net2 VSS INV_D1
x3[3] VDD VOUT net1 VSS INV_D1
x3[2] VDD VOUT net1 VSS INV_D1
x3[1] VDD VOUT net1 VSS INV_D1
x3[0] VDD VOUT net1 VSS INV_D1
.ends

* expanding   symbol:  INV_D1.sym # of pins=4
** sym_path: /home/designer/shared/GRO-TDC/std_cells/INV_D1.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/INV_D1.sch
.subckt INV_D1 VDD VOUT VIN VSS
*.PININFO VDD:B VSS:B VOUT:O VIN:I
M2 VOUT VIN VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

