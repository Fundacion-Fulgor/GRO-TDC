* Extracted by KLayout with SG13G2 LVS runset on : 24/01/2026 20:08

.SUBCKT INV_D1 VIN
M$1 \$1 VIN \$3 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 \$2 VIN \$3 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS INV_D1
