* Extracted by KLayout with SG13G2 LVS runset on : 26/01/2026 15:06

.SUBCKT OR VB VA VSS VDD VOUT
X$1 VSS VDD VA VB \$7 NOR
M$1 VSS \$7 VOUT VSS sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$2 VDD \$7 VOUT VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p PS=1.28u
+ PD=1.28u
.ENDS OR

.SUBCKT NOR \$1 \$2 \$3 VB \$5
M$1 \$5 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.45u AS=0.153p AD=0.153p PS=1.58u
+ PD=1.58u
M$2 \$1 VB \$5 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$3 \$7 \$3 \$2 \$2 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$4 \$5 VB \$7 \$2 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS NOR
