** sch_path: /home/designer/shared/GRO-TDC/GRO.sch
.subckt GRO VDD EN K0 K1 VSS K2
*.PININFO EN:I VDD:B VSS:B K0:O K1:O K2:O
x2 S K0 K2 VSS INV3
x3 S K1 K0 VSS INV3
x4 S K2 K1 VSS INV3
M1 S G VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=32
x5[1]  VDD EN_N EN VSS INV_D1
x5[0]  VDD EN_N EN VSS INV_D1
x6[3]  VDD net1 EN_N VSS INV_D1
x6[2]  VDD net1 EN_N VSS INV_D1
x6[1]  VDD net1 EN_N VSS INV_D1
x6[0]  VDD net1 EN_N VSS INV_D1
x7[7]  VDD net2 net1 VSS INV_D1
x7[6]  VDD net2 net1 VSS INV_D1
x7[5]  VDD net2 net1 VSS INV_D1
x7[4]  VDD net2 net1 VSS INV_D1
x7[3]  VDD net2 net1 VSS INV_D1
x7[2]  VDD net2 net1 VSS INV_D1
x7[1]  VDD net2 net1 VSS INV_D1
x7[0]  VDD net2 net1 VSS INV_D1
x8[15] VDD G net2 VSS INV_D1
x8[14] VDD G net2 VSS INV_D1
x8[13] VDD G net2 VSS INV_D1
x8[12] VDD G net2 VSS INV_D1
x8[11] VDD G net2 VSS INV_D1
x8[10] VDD G net2 VSS INV_D1
x8[9] VDD G net2 VSS INV_D1
x8[8] VDD G net2 VSS INV_D1
x8[7] VDD G net2 VSS INV_D1
x8[6] VDD G net2 VSS INV_D1
x8[5] VDD G net2 VSS INV_D1
x8[4] VDD G net2 VSS INV_D1
x8[3] VDD G net2 VSS INV_D1
x8[2] VDD G net2 VSS INV_D1
x8[1] VDD G net2 VSS INV_D1
x8[0] VDD G net2 VSS INV_D1
M2 S G VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M3 K2 G VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M4 K0 EN_N VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=32
.ends

* expanding   symbol:  /home/designer/shared/GRO-TDC/std_cells/INV3.sym # of pins=4
** sym_path: /home/designer/shared/GRO-TDC/std_cells/INV3.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/INV3.sch
.subckt INV3 VDD VOUT VIN VSS
*.PININFO VDD:B VSS:B VOUT:O VIN:I
x2 VDD net2 VIN VSS INV_D1
x1[1] VDD net1 net2 VSS INV_D1
x1[0] VDD net1 net2 VSS INV_D1
x3[3] VDD VOUT net1 VSS INV_D1
x3[2] VDD VOUT net1 VSS INV_D1
x3[1] VDD VOUT net1 VSS INV_D1
x3[0] VDD VOUT net1 VSS INV_D1
.ends


* expanding   symbol:  /home/designer/shared/GRO-TDC/std_cells/INV_D1.sym # of pins=4
** sym_path: /home/designer/shared/GRO-TDC/std_cells/INV_D1.sym
** sch_path: /home/designer/shared/GRO-TDC/std_cells/INV_D1.sch
.subckt INV_D1 VDD VOUT VIN VSS
*.PININFO VDD:B VSS:B VOUT:O VIN:I
M2 VOUT VIN VDD VDD sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
M1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends

